library verilog;
use verilog.vl_types.all;
entity tb_S_ser is
    generic(
        Clock_Parameter : integer := 64
    );
end tb_S_ser;
