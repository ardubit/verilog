library verilog;
use verilog.vl_types.all;
entity pack_unpack is
end pack_unpack;
