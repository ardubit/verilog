library verilog;
use verilog.vl_types.all;
entity testbench_lab2 is
end testbench_lab2;
