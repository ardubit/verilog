library verilog;
use verilog.vl_types.all;
entity tb is
    generic(
        Clock_Parameter : integer := 64
    );
end tb;
