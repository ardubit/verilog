library verilog;
use verilog.vl_types.all;
entity testbench_lab1 is
end testbench_lab1;
